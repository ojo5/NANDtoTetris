module NOT(
    input wire A,
    output wire X
);
    assign X = ~A;  // Invert A
endmodule

